`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/11/25 15:01:47
// Design Name: 
// Module Name: _2421_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module _2421_tb;
reg clk,rst;
wire z,q3,q2,q1,q0;
_2421 u_2421(clk,rst,z,q3,q2,q1,q0);

initial begin
    clk=1'b1;
    rst=1'b1;
    #30 rst=~rst;
end
always #25 clk=~clk;
initial begin
    #1000
    $finish;
end
endmodule